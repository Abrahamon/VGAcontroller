`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:32:19 09/07/2016 
// Design Name: 
// Module Name:    color_manager 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module color_manager(
    input [5:0] i_seg,
    input [5:0] i_min,
    output [7:0] o_rgb
    );


endmodule
