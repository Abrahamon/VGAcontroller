`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:41:06 09/06/2016 
// Design Name: 
// Module Name:    color_controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module color_controller(
    input wire pixel_pos_x,
	 input wire pixel_pos_y,
	 input wire B_U, B_D, B_L, B_R,B_C,
	 output wire [7:0]rgb
    );


endmodule
